`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:54:55 02/26/2020 
// Design Name: 
// Module Name:    out 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sigmoid(
					clk,
					in,
					out
    );
	 
	 `include "definitions.v"
	 
	 input clk;
	 
	 input wire signed [weight_width-1:0] in;
	 
	 output reg signed [weight_width-1:0] out;
	 
	 reg signed [weight_width-1:0] min_lim = 16'b1111111101000000;
	 reg signed [weight_width-1:0] max_lim = 16'b0000000011000000;
	 
	 always @(posedge clk)
	 begin
		
		if (in < min_lim)
		begin
			out <= 16'b0000000000000000;
		end
		else if (in > max_lim)
		begin
			out <= 16'b0000000000100000;
		end
		else
		begin
			case(in)
				16'b1111111101000000: out <= 16'b0000000000000000;
				16'b1111111101001101: out <= 16'b0000000000000000;
				16'b1111111101011010: out <= 16'b0000000000000000;
				16'b1111111101100110: out <= 16'b0000000000000000;
				16'b1111111101110011: out <= 16'b0000000000000000;
				16'b1111111110000000: out <= 16'b0000000000000001;
				16'b1111111110001101: out <= 16'b0000000000000001;
				16'b1111111110011010: out <= 16'b0000000000000001;
				16'b1111111110100110: out <= 16'b0000000000000010;
				16'b1111111110110011: out <= 16'b0000000000000011;
				16'b1111111111000000: out <= 16'b0000000000000100;
				16'b1111111111001101: out <= 16'b0000000000000101;
				16'b1111111111011010: out <= 16'b0000000000000111;
				16'b1111111111100110: out <= 16'b0000000000001010;
				16'b1111111111110011: out <= 16'b0000000000001101;
				16'b0000000000000000: out <= 16'b0000000000010000;
				16'b0000000000001101: out <= 16'b0000000000010011;
				16'b0000000000011010: out <= 16'b0000000000010110;
				16'b0000000000100110: out <= 16'b0000000000011001;
				16'b0000000000110011: out <= 16'b0000000000011011;
				16'b0000000001000000: out <= 16'b0000000000011100;
				16'b0000000001001101: out <= 16'b0000000000011101;
				16'b0000000001011010: out <= 16'b0000000000011110;
				16'b0000000001100110: out <= 16'b0000000000011111;
				16'b0000000001110011: out <= 16'b0000000000011111;
				16'b0000000010000000: out <= 16'b0000000000011111;
				16'b0000000010001101: out <= 16'b0000000000100000;
				16'b0000000010011010: out <= 16'b0000000000100000;
				16'b0000000010100110: out <= 16'b0000000000100000;
				16'b0000000010110011: out <= 16'b0000000000100000;
				16'b0000000011000000: out <= 16'b0000000000100000;
			endcase
		end
	 end

endmodule
